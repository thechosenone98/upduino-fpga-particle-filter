module particle_filter #(
    parameter string START_MESSAGE = "START_PARTUPDATE",
    parameter string START_MAP_MESSAGE = "START_MAPUPDATE",
) (
    input serial_in,
    output serial_out,
    input clk,
    input reset,
);
    
    wire start_of_particle_message

endmodule